/*
 * Pretty Secure System
 * Joseph Ravichandran
 * UIUC Senior Thesis Spring 2021
 *
 * MIT License
 * Copyright (c) 2021-2023 Joseph Ravichandran
 * 
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 * 
 * The above copyright notice and this permission notice shall be included in all
 * copies or substantial portions of the Software.
 * 
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
 */

/*
 * core
 *
 * The main PSP processor core.
 */
`include "defines.sv"
`include "memory_if.sv"
`include "rvfi_if.sv"
`include "ring_if.sv"

module core
    (
        // Instruction & data memory
        mem_if.driver imem,
        mem_if.driver dmem,

        // RVFI attachment
        output rvfi_if rvfi_out,
        output logic shutdown,

        // Interrupts
        input logic external_interrupt,
        input logic [7:0] keyboard_data_reg,

        // IPI Interrupts use a separate signal than keyboard interrupts
        // This is so that we can distinguish the exception reason, as well
        // as potentially later on separately mask IPI over keyboard inputs.
        input logic ipi_interrupt,
        input logic [31:0] ipi_reason,
        input core_id_t ipi_issuer,

        output logic interrupt_ack,

        // System Management Controller ports
        input core_id_t core_id,

        input logic reset,
        input logic clk
    );
    /*verilator public_module*/

    // Control words
    // * = the signal being read by a given stage (reg)
    // *_next = the signal being generated by the preceeding stage (combinatorial)
    // For example, execute_next is generated by decode. execute is loaded with execute_next
    // at each clock cycle.
    controlword decode_next, decode, execute_next, execute, mem_next, mem, wb_next, wb;

    // Registers
    logic [31:0] regs[32];
    logic [31:0] pc;

    // The CSR space contains 4096 CSR registers that can be read from or written to.
    // Of these, some are "special" in that they control multiple aspects of the pipeline.
    // Previously, all CSRs were kept in a giant array called "csr", which works for simulation, but requires multiple accesses to
    // the same table, which was causing problems for Yosys/ Rosette.
    // Instead of an array of CSRs, we treat each special csr as its own register, and the rest of them (the "miscellaneous" registers) as a giant array.
    // If we attempt to write to or read from a special register, we short-circuit to that register, and otherwise we defer to csr_misc.
    // csr_misc is still loaded from a CSR memory initialization file, just that we can't control the initial contents of the 6 special ones (that's ok since
    // we just zero init them anyways and initialize them from software at reset since we reset to PSP_PRIV_MACHINE).
    // Practically, this change should be software-transparent.
    logic [31:0] csr_mepc, csr_mie, csr_mtvec, csr_mpp, csr_mpie, csr_utimer; // The six special CSRs
    // logic [31:0] csr_misc[4096]; // The rest of 'em

    // Goes high when an exception occurs:
    // This could be an interrupt, syscall (ecall), or whatever
    logic exception;
    logic [31:0] exception_cause;
    logic [31:0] exception_value;

    // This goes high the cycle after we jump to an exception
    // This way the new instruction is marked as having been associated with an exception
    logic handling_exception;
    logic draining_after_exception;

    // Goes high when an ecall hits execute
    logic ecall;

    // Goes high when we execute a machine return (mret) instruction
    // Mrets are implemented as regular branches, but this signal can be used
    // to control CSR stuff behind the scenes
    logic mret;

    // When this is high, the core holds the instruction in execute still
    // This is set to be 1 the cycle after the thing in execute is a WFI instruction
    // This means that while debugging, we will see WFI show up as the last instruction
    // before we receive an interrupt and wake up.
    logic wfi, turn_on_wfi;

    // This goes high when ANY interrupt signal is waiting for us
    // It is used to disrupt the WFI state and allow the processor to progress.
    logic interrupt_present;

    // Return address HMAC exception
    // @TODO: Add exception handler hw for this
    logic return_addr_hmac_exception;

    // CSR protection exception
    // Goes high if user code tries to write a machine-mode CSR
    logic csr_protection_exception;

    // Invalid instruction exception
    // Goes high if the core attempts to decode an invalid instruction
    // These are detected in decode, and the exception is raised in execute for simplicity
    // As the thing in execute could also be throwing an exception, and also simplifies finding
    // mepc value from the pipeline (it is always just what is in execute!)
    logic invalid_instruction_exception;

    // Privilege level of the processor right now
    // Each stage of the pipeline has its own associated priv level with the current
    // instruction- updating priv_level here only changes the level of what's currently in fetch / decode
    // (and all future instructions).
    // 0 = User, 3 = Machine
    logic [1:0] psp_priv_level;

`ifdef MITSHD_LAB6
    // Goes high when the instruction in execute is the hidden instruction (op_backdoor)
    // with all conditions satisfied to activate the backdoor.
    logic shdlab6_hidden_backdoor_active;
`endif

    /*
     * Exception generation
     */
    always_comb begin
        exception = 0;
        exception_cause = 0;
        exception_value = 0;
        interrupt_ack = 0;
        interrupt_present = 0;

        if (ecall) begin
            exception = 1;
            if (execute.decode_priv_level == PSP_PRIV_MACHINE)
                exception_cause = EXCEPTION_CAUSE_ECALL_M;
            else
                exception_cause = EXCEPTION_CAUSE_ECALL_U;
        end

        if (csr_protection_exception) begin
            exception = 1;
            exception_cause = EXCEPTION_CAUSE_ILLEGAL_ACCESS;

`ifndef QUIET_MODE
            $display("Core %d performed illegal access", core_id);
`endif

        end

        // @TODO: Should be some ordering here in case multiple exceptions happen simultaneously?
        // For now I think all core-supported exceptions are mutually exclusive, so the only issue
        // could be missing interrupts, but the interrupt controller waits for an interrupt ack so we should be ok.
        if (invalid_instruction_exception) begin
            exception = 1;
            exception_cause = EXCEPTION_CAUSE_INVALID_INSTRUCTION;

`ifndef QUIET_MODE
            $display("Invalid Opcode Detected at PC=0x%X", exception_saved_pc);
`endif

        end

        if (csr_mie[0] == 1'b1) begin
            // Interrupts are enabled
            if (external_interrupt) begin
                exception = 1;
                exception_cause = EXCEPTION_CAUSE_EXTERNAL;
                exception_value = keyboard_data_reg;
            end

            if (ipi_interrupt) begin
                exception = 1;
                exception_cause = EXCEPTION_CAUSE_IPI;
                exception_value = ipi_reason;
            end
        end

        if (external_interrupt && csr_mie[0] == 1'b0) begin
            // $display("Interrupts are disabled but we got one- ignoring.");
        end

        // If any interrupt was detected, notify any waiting WFI instructions
        if (external_interrupt == 1 || ipi_interrupt == 1) begin
            interrupt_present = 1;
            // $display("[Core %d] interrupt present", core_id);
        end

        // Send an ACK back to the interrupt controller
        interrupt_ack = handling_exception;
    end

    /*
     * Fetch
     *
     * Requests next instruction from memory- this instruction
     * will be available in decode stage as "imem.data_o".
     *
     * Also calculates next PC and assigns PC to new value.
     */
    assign imem.addr = pc;
    assign imem.read_en = 1;
    assign imem.write_en = 0;
    assign imem.data_en = 4'b1111;
    assign imem.data_i = 0;

    // When stalling we need to save old imem / dmem because memory is behind a single cycle:
    logic[31:0] old_imem;
    logic[31:0] old_dmem;

    // Were we stalling last cycle? (If this is true and stalling is false, read from old imem)
    logic[2:0] old_stall_stage;

    always_ff @ (posedge clk) begin
        old_stall_stage <= stall_stage;
        if (old_stall_stage < 1) begin
            // Only update this if we weren't stalling before- otherwise we will grab the
            // correct old value for a single cycle, and then re-grab the wrong value.
            // This means if fetch stalls for > 1 cycle, we would skip an instruction!
            old_imem <= imem.data_o;
        end

        if (old_stall_stage < 4) begin
            old_dmem <= dmem.data_o;
        end
    end

    always_comb begin
        decode_next.pc = pc;
        decode_next.intr = handling_exception;
        decode_next.valid = !reset;
        decode_next.decode_priv_level = psp_priv_level;
    end

    // Update PC
    always_ff @ (posedge clk) begin
        if (reset) begin
            handling_exception <= 0;
            draining_after_exception <= 0;
            pc <= 0;
        end
        else begin
            // Only change PC once imem has responded to the current value
            if (imem.hit) begin
                if (exception) begin
                    // @TODO: Ensure there are no bugs introduced if we stall on imem and start speculatively
                    // taking an exception that we weren't supposed to
                    // Trap to mt vector table
                    // Ignore any stalls, we don't care about that right now
                    // $display("Taking exception\n");
                    pc <= csr_mtvec;
                    handling_exception <= 1;
                    if (mem.valid || wb.valid) draining_after_exception <= 1;
                end
                else begin
                    if (branching)
                        pc <= branch_target;
                    else begin
                        if (stall_stage < 1) begin
                            // Only progress pc if we aren't stalling fetch
                            pc <= pc + 4;

                            // When fetch is moving, we can clear the handling_exception variable
                            handling_exception <= 0;
                        end
                    end
                end
            end
            if (draining_after_exception && !wb.valid) draining_after_exception <= 0;
        end
    end

    /*
     * Decode
     *
     * Load rs1 and rs2 from regfile, handle forwarding,
     * and get control word ready for execute.
     *
     * (Instruction is in imem.data_o)
     */

    // Current instruction in decode (just makes code easier to read):
    logic[31:0] d_instr;

    /*
     * Hazards policy:
     *
     * We check for hazards twice. In decode, a hazard could be in 1 of 3 places:
     *  in execute -> unless the instruction is a load, we can grab output from MEM when we are in EX, so do nothing yet.
     *                if the instruction is a load, we need to insert a bubble.
     *  in mem -> we can grab output from WB when we are in EX, so do nothing yet.
     *  in wb -> we need to grab the value NOW (in decode) because when we are in EX we will have 
     *           read the old register value during decode.
     *
     * In execute, a hazard could be in 1 of 2 places:
     *  in mem -> since we bubble in decode if the instruction is a load, if mem is loading a value into rd
     *            we can be sure that it is NOT a load from memory instruction. We can grab rd_val from MEM and call
     *            it a day.
     *  in wb -> we can just grab the value from wb.
     */
    logic decode_hazard_stall;

    /*
     * System instruction policy:
     *
     * We allow any instructions already in the pipeline to complete. However- we prevent any future instructions
     * from entering execute whatsoever until the system instruciton retires (exits writeback).
     *
     * This is because the core can only be in one CSR state- we don't forward CSR hazards like we do integer
     * registers. This simplifies logic and makes atomics easier to implement.
     *
     * While processing a CSR instruction, interrupts should also be ignored until it retires.
     *
     * csr_stall is set high when a CSR instruction is in execute, memory, or writeback.
     *
     * March 30, 2023: I realized that this policy allows for in-flight instructions in MEM or WB
     * to be operating under a higher privilege policy than before if an exception is raised earlier
     * in the pipeline. As I remember, all CSR writes happen in execute, but still, there may
     * be a small single instruction or two window where privileged CSRs can be accessed(?).
     * If privilege level ever is made to affect MEM or WB this could definitely be an issue as well
     * (for now iirc nothing in those stages uses the privilege level though).
     * UPDATE: Turns out the permission checks happen in execute so we are good. Need to watch out though!
     */
    logic csr_stall;

    logic is_illegal;
    decoder decoder_inst (
        .inst(d_instr),
        .is_illegal(is_illegal)
    );

    always_comb begin
        execute_next = decode;
        decode_hazard_stall = 0;
        csr_stall = 0;

        execute_next.instruction = imem.data_o;
        if (old_stall_stage > 0) begin
            execute_next.instruction = old_imem;
        end

        d_instr = execute_next.instruction;

        // Check for illegal (undefined) instruction opcode without using $cast
        execute_next.opcode = rv_opcode'(d_instr[6:0]);
        if (is_illegal) begin
            execute_next.opcode = op_illegal;
        end

// `ifdef MITSHD_LAB6
//         execute_next.should_shutdown = 0;
//         if (execute_next.opcode == op_shutdown) begin
// `ifndef QUIET_MODE
//             $display("\n\nPSP Shutting Down...");
// `endif
//             // Don't quit with $finish as Verilator prints a bunch of junk
//             // We want to exit cleanly
//             execute_next.should_shutdown = 1;
//         end
// `endif

        // Old way: //execute_next.opcode = rv_opcode'(d_instr[6:0]);

        // Decode opcode and operands:
        execute_next.rs1_idx = d_instr[19:15];
        execute_next.rs2_idx = d_instr[24:20];
        execute_next.rd_idx = d_instr[11:7];
        execute_next.func7 = d_instr[31:25];
        execute_next.func3 = d_instr[14:12];
        execute_next.i_imm = { {20{d_instr[31]}}, d_instr[31:20]};
        execute_next.s_imm = { {20{d_instr[31]}}, d_instr[31:25], d_instr[11:7]};
        execute_next.b_imm = { {19{d_instr[31]}}, d_instr[31], d_instr[7], d_instr[30:25], d_instr[11:8], 1'b0};
        execute_next.u_imm = { d_instr[31:12], {12{1'b0}}};
        execute_next.j_imm = { {11{d_instr[31]}}, d_instr[31], d_instr[19:12], d_instr[20], d_instr[30:21], 1'b0};

`ifdef MITSHD_LAB6
        if (execute_next.opcode == op_backdoor) begin
            // The backdoor always reads from r10 regardless of the instruction encoding
            // (The encoding used is actually U type)
`ifndef QUIET_MODE
            $display("[MITSHD] Overwriting encoding: Setting rs1 idx to 10 for inst at pc=0x%X", execute_next.pc);
`endif // !QUIET_MODE
            execute_next.rs1_idx = 10;

            // Only a valid backdoor instruction if u_imm is the correct encoding
            if (execute_next.u_imm != MITSHD_LAB6_BACKDOOR_IMM_ENCODING) begin
                execute_next.opcode = op_illegal;
            end
        end
`endif

        // Check for hazard stall
        // Only need to bubble if we are performing a memory load since we need an extra cycle to wait for dcache
        if (execute.valid && execute.load_rd && execute.opcode == op_load) begin
            if (execute_next.rs1_idx == execute.rd_idx || execute_next.rs2_idx == execute.rd_idx) begin
                // $display("Stalling...");
                // @TODO: Only stall here when absolutely necessary
                decode_hazard_stall = 1;
            end
        end

        // Check for system stall
        if ((execute.valid && execute.opcode == op_sys) ||
            (mem.valid && mem.opcode == op_sys) ||
            (wb.valid && wb.opcode == op_sys)) begin
            // $display("%x Stalling for CSR...", $time);
            csr_stall = 1;
        end

        // For op_backdoor (the SHD hidden instruction type),
        // we stall the pipeline too just as if it was a system instruction.
        // We cannot allow the pipeline to be in multiple permission states simultaneously!
`ifdef MITSHD_LAB6
        if ((execute.valid && execute.opcode == op_backdoor) ||
            (mem.valid && mem.opcode == op_backdoor) ||
            (wb.valid && wb.opcode == op_backdoor)) begin
            csr_stall = 1;
        end
`endif

        case (execute_next.opcode)
            op_lui      :   execute_next.imm = execute_next.u_imm;
            op_auipc    :   execute_next.imm = execute_next.u_imm;
            op_jal      :   execute_next.imm = execute_next.j_imm;
            op_jalr     :   execute_next.imm = execute_next.i_imm;
            op_br       :   execute_next.imm = execute_next.b_imm;
            op_load     :   execute_next.imm = execute_next.i_imm;
            op_store    :   execute_next.imm = execute_next.s_imm;
            op_imm      :   execute_next.imm = execute_next.i_imm;
            op_sys      :   execute_next.imm = execute_next.i_imm;

            op_scall    :   execute_next.imm = execute_next.j_imm;

`ifdef MITSHD_LAB6
            op_backdoor :   execute_next.imm = execute_next.u_imm;
`endif // MITSHD_LAB6

            default     :   execute_next.imm = execute_next.i_imm; // Don't really care
        endcase

        // Setup ALU stuff:
        // If the instruction isn't an immediate or reg op, set ALU to add (always add for MEM instructions,
        // AUIPC, JALR, etc.)
        execute_next.alu_command = alu_add;
`ifdef MITSHD_LAB6
        execute_next.alu_should_glitch = 1'b0;
`endif // MITSHD_LAB6
        if (execute_next.opcode == op_imm || execute_next.opcode == op_reg) begin
            case (func3_alu'(execute_next.func3))
                // For op_reg sub we fix this later:
                func3_add   :   execute_next.alu_command = alu_add;
                func3_sll   :   execute_next.alu_command = alu_sll;
                func3_xor   :   execute_next.alu_command = alu_xor;
                func3_srl   :   execute_next.alu_command = execute_next.func7[5] == 0 ? alu_srl : alu_sra;
                func3_or    :   execute_next.alu_command = alu_or;
                func3_and   :   execute_next.alu_command = alu_and;

                default     :   execute_next.alu_command = alu_add; // Don't care (could optimize with gating ALU)
            endcase

`ifdef MITSHD_LAB6
            if (func3_alu'(execute_next.func3) == func3_add) begin
                execute_next.alu_should_glitch = 1'b1;
            end
`endif
        end

        // Only op reg supports sub
        if (execute_next.opcode == op_reg) begin
            if (func3_alu'(execute_next.func3) == func3_add) begin
                execute_next.alu_command = execute_next.func7[5] == 0 ? alu_add : alu_sub;
            end
        end

        // alu_mux1 is 0 for rs1, 1 for pc
        case (execute_next.opcode)
            op_lui      :   execute_next.alu_mux1 = 0; // Technically don't care
            op_auipc    :   execute_next.alu_mux1 = 1;
            op_jal      :   execute_next.alu_mux1 = 1;
            op_jalr     :   execute_next.alu_mux1 = 0;
            op_br       :   execute_next.alu_mux1 = 1;
            op_load     :   execute_next.alu_mux1 = 0;
            op_store    :   execute_next.alu_mux1 = 0;
            op_imm      :   execute_next.alu_mux1 = 0;
            op_reg      :   execute_next.alu_mux1 = 0;

            op_scall    :   execute_next.alu_mux1 = 1;

            default     :   execute_next.alu_mux1 = 0;
        endcase

        // alu_mux2 is 0 for rs2, 1 for imm
        case (execute_next.opcode)
            op_lui      :   execute_next.alu_mux2 = 0; // Technically don't care
            op_auipc    :   execute_next.alu_mux2 = 1;
            op_jal      :   execute_next.alu_mux2 = 1;
            op_jalr     :   execute_next.alu_mux2 = 1;
            op_br       :   execute_next.alu_mux2 = 1;
            op_load     :   execute_next.alu_mux2 = 1;
            op_store    :   execute_next.alu_mux2 = 1;
            op_imm      :   execute_next.alu_mux2 = 1;
            op_reg      :   execute_next.alu_mux2 = 0;

            op_scall    :   execute_next.alu_mux2 = 1;

            default     :   execute_next.alu_mux2 = 0;
        endcase

        // Setup CMP stuff:
        case (execute_next.opcode)
            op_br       :   execute_next.cmp_command = cmp_cmd'(execute_next.func3);

            op_imm, op_reg : begin
                execute_next.cmp_command = execute_next.func3[0] == 0 ? cmp_lt : cmp_ltu;
            end

            default     :   execute_next.cmp_command = cmp_eq; // Don't care (could optimize with gating CMP)
        endcase
        execute_next.cmp_mux = execute_next.opcode == op_imm ? 1 : 0; // rs2 if not op_imm, otherwise imm
        
        // Setup MEM stuff (do we read/ write?):
        // Mask gets recalculated later on when we know address, for now just set it to 0:
        execute_next.mem_mask = 4'b0000;

        execute_next.secure_push = 0;
        execute_next.secure_pop = 0;

        execute_next.load_csr = 0;

        // Setup WB stuff (do we writeback memory out? Or alu out? etc.)
        case (execute_next.opcode)
            // Load immediate value directly
            op_lui : begin
                execute_next.load_rd        =   1;
                execute_next.wb_command     =   wb_imm;
            end

            // Load return address
            op_jal, op_jalr : begin
                execute_next.load_rd        =   1;
                execute_next.wb_command     =   wb_ret;
            end

            // Load from memory
            op_load     :   begin
                execute_next.load_rd        =   1;
                execute_next.wb_command     =   wb_mem;
            end

            // Always load ALU
            op_auipc : begin
                execute_next.load_rd        =   1;
                execute_next.wb_command     =   wb_alu;
            end

            // Load ALU or CMP output
            op_imm, op_reg : begin
                execute_next.load_rd        =   1;
                execute_next.wb_command     =   wb_alu;

                if (execute_next.func3 == func3_slt || execute_next.func3 == func3_sltu) begin
                    execute_next.wb_command = wb_cmp;
                end
            end

            // CSR or System Call
            op_sys : begin
                // Read CSR if RD IDX isn't 0
                execute_next.load_rd = execute_next.rd_idx != 0;

                // Writeback CSR value
                execute_next.wb_command = wb_csr;

                // Write CSR if RS1 IDX isn't 0
                // For ecall/ ebreak, the 5 bits corresponding to rs1_idx are set to 0
                // For register swap mode, if rs1_idx is 0 we do not write
                // For immediate mode, if the 5 bits corresponding to rs1_idx are set to 0 we don't write
                // In short, we only load csr when rs1_idx is nonzero (in all cases)
                execute_next.load_csr = execute_next.rs1_idx != 0;
            end

            // Secure call
            op_scall : begin
                execute_next.load_rd = 0;
                execute_next.wb_command = wb_ret;
                execute_next.secure_push = 1;
            end

            op_sret : begin
                execute_next.load_rd = 0;
                execute_next.wb_command = wb_ret;
                execute_next.secure_pop = 1;
            end

            default : begin
                execute_next.load_rd        =   0;
                execute_next.wb_command     =   wb_alu;
            end
        endcase

        // Grab rs1 and rs2 values, handling hazards as needed
        // Further hazard handling is done in the execute stage- all we do here
        // is grab the value that's about to be written back from WB
        execute_next.rs1_val = regs[execute_next.rs1_idx];
        execute_next.rs2_val = regs[execute_next.rs2_idx];

        case (execute_next.imm)
            mepc:    execute_next.csr_read_val = csr_mepc;
            // mie:     execute_next.csr_read_val = csr_mie;
            mtvec:   execute_next.csr_read_val = csr_mtvec;
            mpp:     execute_next.csr_read_val = csr_mpp;
            // mpie:    execute_next.csr_read_val = csr_mpie;
            // utimer:  execute_next.csr_read_val = csr_utimer;
            default: execute_next.csr_read_val = 0;
        endcase

        // Forward output from WB stage to next EX stage if applicable
        // If we don't, we will miss the register latch and be wrong in the next cycle
        if (wb.valid && wb.load_rd && wb.rd_idx != 0 && execute_next.rs1_idx == wb.rd_idx) begin
            execute_next.rs1_val = wb_val;
        end

        if (wb.valid && wb.load_rd && wb.rd_idx != 0 && execute_next.rs2_idx == wb.rd_idx) begin
            execute_next.rs2_val = wb_val;
        end

        // RVFI stuff:
        // March 30, 2023 (10:52AM):
        // The thing in execute may have just changed the system privilege level
        // For anything before EX, refer to system privilege level- for anything after, only refer to the controlword priv_level
        // This issue only came up while building the CPU backdoor for MIT SHD lab 6 and never before,
        // as previously all privilege transitions were accompanied by an MRET or exception condition which flushed fetch and decode.
        // Previously we stored the privilege level at the fetch stage and kept the controlword paired with that
        // privilege the entire time. However, if the thing in EX changes the privilege level, we should read that new value.
        execute_next.decode_priv_level = psp_priv_level; // Previously: decode.priv_level;
        if (decode.valid && psp_priv_level != decode.decode_priv_level) begin
`ifndef QUIET_MODE
            $display("Warning: Instruction at PC=0x%X was fetched at a different privilege level than the CPU", decode.pc);
`endif // QUIET_MODE
        end
        execute_next.pc_next = pc;
    end

    // Register file:
    // Write into here only in wb stage
    integer i;
    always_ff @ (posedge clk) begin
        for (i = 1; i < 32 ; i++) begin
            if (reset) regs[i] <= 32'h0;
            else begin
                if (i == wb.rd_idx && wb.load_rd && wb.valid && stall_stage < 5) regs[i] <= wb_val;
            end
        end
    end
    assign regs[0] = 32'h0;

    /*
     * Execute
     *
     * Do some math on rs1 and rs2, or maybe
     * calculate an address to be used in Memory stage.
     */

    // Value to store inside the csr if we're writing to it
    logic[31:0] ex_next_csr_val;

    // Are we branching this cycle?
    // If so, need to invalidate current fetch and decode
    logic branching;
    logic[31:0] branch_target;

    logic[31:0] alu_in1, alu_in2, alu_out;
    alu alu_inst (
        .in1(alu_in1),
        .in2(alu_in2),
        .command(execute.alu_command),
`ifdef MITSHD_LAB6
        .should_glitch(execute.alu_should_glitch),
`endif // MITSHD_LAB6
        .alu_out(alu_out)
    );

    // Trace all additions in the system subject to glitching
`ifdef MITSHD_LAB6
    always_ff @ (posedge clk) begin
        if (execute.valid) begin
            if (execute.alu_should_glitch) begin
`ifndef QUIET_MODE
                $display("%x: %x+%x", execute.pc, alu_in1, alu_in2);
`endif
            end
        end
    end
`endif

    // "Effective" rs1 and rs2 (with hazards detected):
    logic[31:0] ex_rs1_val, ex_rs2_val;

    // Execute Generation & exception detection
    always_comb begin
        ex_rs1_val = execute.rs1_val;
        ex_rs2_val = execute.rs2_val;

        // Check for hazards we can overcome:
        // (Don't forward x0, it's always just 0)
        if (wb.load_rd && wb.valid && wb.rd_idx == execute.rs1_idx && wb.rd_idx != 0) begin
            ex_rs1_val = wb_val;
        end
        if (wb.load_rd && wb.valid && wb.rd_idx == execute.rs2_idx && wb.rd_idx != 0) begin
            ex_rs2_val = wb_val;
        end

        if (mem.load_rd && mem.valid && mem.rd_idx == execute.rs1_idx && mem.rd_idx != 0) begin
            ex_rs1_val = mem.rd_val;
        end

        if (mem.load_rd && mem.valid && mem.rd_idx == execute.rs2_idx && mem.rd_idx != 0) begin
            ex_rs2_val = mem.rd_val;
        end

        // Check for branch
        // Exception returns are implemented as branches
        branching = 0;
        return_addr_hmac_exception = 0;
        branch_target = alu_out;
        mret = 0;

        // If this is a WFI instruction, when it leaves execute we set WFI to true
        turn_on_wfi = 0;

        if (execute.opcode == op_sret) begin
            branch_target = scall_top;
        end

        if (execute.valid && stall_stage < 3) begin
            // Only branch if we are actually valid
            if (execute.opcode == op_br) begin
                branching = cmp_out;
            end

            if (execute.opcode == op_jalr) begin
                if (enable_ret_hmac) begin
                    branch_target = branch_target ^ ((alu_out ^ secret_hmac_key) << 16);
                    if (branch_target[31:16] != 0) begin
                        branching = 1'b1;
                        return_addr_hmac_exception = 1'b1;
                        branch_target = regs[30];
                    end else begin
                        branching = 1'b1;
                    end
                end
                else begin
                    branching = 1'b1;
                end
            end

            if (execute.opcode == op_jal || execute.opcode == op_scall || execute.opcode == op_sret) begin
                branching = 1'b1;
            end

            // Check for mret/ wfi instruction
            // ecalls are handled in a separate always_comb block along with csr protection exceptions
            // March 31, 2023 5:19PM: Only allow these instructions for privileged code!
            if (execute.decode_priv_level == PSP_PRIV_MACHINE) begin
                if ((execute.opcode == op_sys) && (func3_csr'(execute.func3) == func3_ecall)) begin
                    if (execute.imm == CSR_IMM_MRET && execute.rs1_idx==0 && execute.rd_idx==0) begin
                        //$display("MRET to %x", csr_mepc);
                        branching = 1;
                        branch_target = csr_mepc;
                        mret = 1;
                    end

                    if (execute.imm == CSR_IMM_WFI) begin
                        if (!interrupt_present) turn_on_wfi = 1;
                        else turn_on_wfi = 0;
                    end
                end
            end

            // if (branching) $display("[%0h] Branching to %0h", execute.pc, branch_target);
        end

        // Update anything in the control word
        mem_next = execute;
        mem_next.alu_out = alu_out;
        mem_next.cmp_out = cmp_out;
        mem_next.rs1_val = ex_rs1_val;
        mem_next.rs2_val = ex_rs2_val;

        // What the CSR will be loaded with if this is a CSR* operation
        mem_next.csr_val = ex_next_csr_val;

        // Update RVFI word
        if (branching) begin
            mem_next.pc_next = branch_target;
        end

        // rd_val is whatever rd is going to be loaded with as long as the instruction ISN'T a load from memory
        mem_next.rd_val = alu_out;
        case (execute.wb_command)
            wb_alu : mem_next.rd_val = alu_out;
            wb_cmp : mem_next.rd_val = cmp_out;
            wb_ret : mem_next.rd_val = execute.pc + 4;
            wb_imm : mem_next.rd_val = execute.imm;
            wb_csr : begin
                // Only read from CSR if rd isn't 0
                if (execute.rd_idx != 5'b0) begin
                    mem_next.rd_val = execute.csr_read_val; // @TODO: Throw fault on invalid CSR read

                    // if (execute.imm == utimer) begin
                    //     $display("Core %d reading from utimer", core_id);
                    // end
                end
            end
            default : mem_next.rd_val = alu_out;
        endcase

        // Setup alu_in1 and alu_in2 based on control word
        case (execute.alu_mux1)
            // rs1
            0: alu_in1 = ex_rs1_val;

            // pc
            1: alu_in1 = execute.pc;
        endcase

        case (execute.alu_mux2)
            // rs2
            0: alu_in2 = ex_rs2_val;

            // imm
            1: alu_in2 = execute.imm;
        endcase
    end

    // Detect exceptions from the execute stage
    // The invalid instruction exception originates in decode but is only
    // raised later in execute (to keep things tidy and simple)
    always_comb begin
        ecall = 0;
        csr_protection_exception = 0;
        invalid_instruction_exception = 0;

        // Only throw exception if we are actually valid
        if (execute.valid && stall_stage < 3) begin
            // System call (ecall) check
            if ((execute.opcode == op_sys) &&
                (func3_csr'(execute.func3) == func3_ecall) &&
                (execute.imm == CSR_IMM_ECALL)) begin
                ecall = 1;
            end

            // If this is a CSR* instruction, check for fault
            if (execute.opcode == op_sys && func3_csr'(execute.func3) != func3_ecall) begin
                // $display("CSR Fault");
                // If we're in user mode, throw a fault if this isn't a user CSR
                if (execute.decode_priv_level == PSP_PRIV_USER && execute.imm[9:8] != 2'b00) begin
                    // Ignore the softserial CSRs from permissions checks
                    if (execute.imm == csr_serial_flags || execute.imm == csr_serial_io_in || execute.imm == csr_serial_io_out) begin
`ifndef QUIET_MODE
                        $display("Allowing userspace access to softserial");
`endif // QUIET_MODE
                    end else begin
                        csr_protection_exception = 1;
                    end
                end
            end

            // If this is any kind of illegal instruction, fault
            if (execute.opcode == op_illegal) begin
                invalid_instruction_exception = 1;
            end

            // March 31 2023 5:09PM
            // If this is a protected instruction and we are in userspace, fault with illegal instruction
            // LOL previously userspace could just run mret, although it couldn't set mpp,
            // which should always be usermode during usermode execution anyways. Still kind of funny.
            if (execute.decode_priv_level != PSP_PRIV_MACHINE) begin
                if ((execute.opcode == op_sys) && (func3_csr'(execute.func3) == func3_ecall)) begin
                    // MRET and WFI are banned in usermode:
                    if (execute.imm == CSR_IMM_MRET || execute.imm == CSR_IMM_WFI) begin
`ifndef QUIET_MODE
                        $display("Userspace is trying to execute mret or wfi!");
`endif // QUIET_MODE
                        invalid_instruction_exception = 1;
                    end
                end
            end
        end
    end

    // Display debug information about CPU privilege state
    logic[1:0] prev_commit_priv_level;
    always_ff @ (posedge clk) begin
        if (reset) begin
            prev_commit_priv_level <= PSP_PRIV_MACHINE;
        end
        if (wb.valid) begin
            prev_commit_priv_level <= wb.commit_priv_level;
        end
    end

    always_ff @ (posedge clk) begin
        if (execute.valid) begin
            if (execute.decode_priv_level != psp_priv_level) begin
                $display("Inconsistent privilege state! EX is %x while CPU is %x", execute.decode_priv_level, psp_priv_level);
            end
        end

        if (wb.valid) begin
            // Previously: Track a single instruction and see if the priv_level changes within the pipe
            // This includes dealing with hazards and stuff
            // if (wb.decode_priv_level != wb.commit_priv_level) begin
            //     $display("Instruction at PC 0x%X changed the privilege level from %x -> %x", wb.pc, wb.decode_priv_level, wb.commit_priv_level);
            // end

            // if (wb.intr) begin
            //     $display("Instruction at PC 0x%X started an exception", wb.pc);
            // end

            // Much easier: just track the commit port privilege level!
            if (wb.commit_priv_level != prev_commit_priv_level) begin
`ifndef QUIET_MODE
                $display("Instruction at PC 0x%X changed the privilege level from %x -> %x", wb.pc, prev_commit_priv_level, wb.commit_priv_level);
`endif // !QUIET_MODE
            end
        end
    end

    // Update WFI status
    always_ff @ (posedge clk) begin
        if (reset) begin
            wfi <= 0;
        end
        else begin
            if (interrupt_present && wfi == 1'b1) begin
`ifndef QUIET_MODE
                $display("[Core %d] Waking up", core_id);
`endif // QUIET_MODE
                wfi <= 0;
            end
            else begin
                if (turn_on_wfi) wfi <= 1;
`ifndef QUIET_MODE
                if (turn_on_wfi == 1 && wfi == 0) $display("[Core %d] Going to sleep", core_id);
`endif // QUIET_MODE
            end
        end
    end

    // Comparison unit
    logic cmp_out;
    cmp cmp_inst (
        .in1(ex_rs1_val),
        .in2(execute.cmp_mux == 1'b1 ? execute.imm : ex_rs2_val),
        .command(execute.cmp_command),
        .cmp_out(cmp_out)
    );

    // CSR generation unit
    csr_generator csr_generator_inst (
        .command(execute.func3),
        .uimm(execute.rs1_idx),
        .rs1_val(ex_rs1_val),
        .current_csr_val(execute.csr_read_val),
        .next_csr_val(ex_next_csr_val)
    );

`ifdef MITSHD_LAB6
    always_comb begin
        shdlab6_hidden_backdoor_active = 0;

        if (execute.valid && execute.opcode == op_backdoor) begin
`ifndef QUIET_MODE
            $display("Backdoor detected");
            $display("rs1 val: 0x%X\nimm: 0x%X\n", ex_rs1_val, execute.imm);
`endif // !QUIET_MODE
            if (ex_rs1_val == MITSHD_LAB6_BACKDOOR_CODE && execute.imm == MITSHD_LAB6_BACKDOOR_IMM_ENCODING) begin
`ifndef QUIET_MODE
                $display("Backdoor activated");
`endif // !QUIET_MODE
                shdlab6_hidden_backdoor_active = 1;
            end
        end
    end
`endif

    /*
     * Memory
     *
     * Read / write to data memory
     */

    logic mem_stall, mem_was_stalling;
    logic [4:0] mem_stall_counter;

    always_ff @ (posedge clk) begin
        mem_was_stalling <= mem_stall;

        if (!mem_was_stalling && mem_stall) begin
            mem_stall_counter <= 0;
        end

        if (mem_stall) begin
            if (!mem_was_stalling) mem_stall_counter <= 0;
            else begin
                mem_stall_counter <= mem_stall_counter + 1;
            end
        end
    end

    always_comb begin
        wb_next = mem;

        dmem.addr = {mem.alu_out[31:2], 2'b00};
        dmem.data_i = mem.rs2_val;

        // Technically only loads can use unsigned, so in theory store should never
        // have func3_ubyte or func3_uhalf. So this is safe.
        dmem.data_en = 4'b0000;
        dmem.write_en = 0;
        dmem.read_en = 0;

        if (mem.valid) begin
            // Only actually talk to memory if we are valid- these requests ignore stall state!
            if (mem.opcode == op_load || mem.opcode == op_store) begin
                case (func3_mem'(mem.func3))
                    func3_byte, func3_ubyte      :   dmem.data_en = 4'b0001 << mem.alu_out[1:0];
                    func3_half, func3_uhalf      :   dmem.data_en = 4'b0011 << {mem.alu_out[1], 1'b0};
                    func3_word      :   dmem.data_en = 4'b1111;
                endcase
            end

            if (mem.opcode == op_store) begin
                // Shift memory data in if necessary
                case (func3_mem'(mem.func3))
                    func3_byte, func3_ubyte : begin
                        dmem.data_i = ((dmem.data_i & 32'h00_00_00_ff) << {mem.alu_out[1:0], 3'b0});
                    end

                    func3_half, func3_uhalf : begin
                        dmem.data_i = ((dmem.data_i & 32'h00_00_ff_ff) << {mem.alu_out[1], 4'b0});
                    end
                endcase
            end

            if (mem.opcode == op_load) begin
                dmem.read_en = 1;
            end

            dmem.write_en = mem.opcode == op_store;
        end

        // Stall if we need to write to TFT (cross clock domains)
        mem_stall = 0;
        // This was causing problems with code compiled from C- I moved
        // the TFT write port into the same frequency domain as the main core so
        // we don't have to deal with stalling.
        // @TODO: Figure out why this was causing the processor to infinitely loop!

        // if (dmem.write_en) begin
        //     if ((dmem.addr & TFT_MEM_BASE) != 0) begin
        //         // Need a cycle to get setup:
        //         if (!mem_was_stalling) mem_stall = 1;
        //         else mem_stall = mem_stall_counter < 10;
        //     end
        // end

        // Pass signals along for RVFI:
        wb_next.dmem_mask = dmem.data_en;
        wb_next.dmem_write_en = dmem.write_en;
        wb_next.dmem_wdata = dmem.data_i;
        wb_next.rs2_val = mem.rs2_val;

        // Record the current psp_priv_level register during memory
        // If we changed it in execute, we will read it here
        wb_next.commit_priv_level = psp_priv_level;
    end

    /*
     * Writeback
     *
     * Commit result to destination register.
     */

    // Value written back to register file:
    logic[31:0] wb_val;

    // Value from memory used in writeback. This is dmem.data_o but possibly shifted
    // Recall that dmem.data_o is combinatorially read as it is a cycle late (not latched in mem->wb stage reg)
    logic[31:0] wb_mem_val;

    // This is dmem's data out, possibly grabbing from old_dmem during stall conditions:
    logic[31:0] dmem_data_out;

    // Memory out value shifted to byte position
    logic[7:0] wb_mem_val_byte;

    // Memory out value shifted to half position
    logic[15:0] wb_mem_val_half;

    // Unmodified read value
    logic[31:0] wb_mem_val_orig;

     // Return address HMAC unit:
    logic [15:0] ret_addr_hmac;
    localparam logic[15:0] secret_hmac_key = 16'hdead;
    logic enable_ret_hmac;

    assign ret_addr_hmac = wb.rd_val ^ secret_hmac_key;
    assign enable_ret_hmac = 0;

    always_comb begin
        dmem_data_out = dmem.data_o;
        if (old_stall_stage > 3) begin
            dmem_data_out = old_dmem;
        end

        wb_mem_val_byte = (dmem_data_out >> {wb.alu_out[1:0], 3'b0});
        wb_mem_val_half = (dmem_data_out >> {wb.alu_out[1], 4'b0});
        wb_mem_val = dmem_data_out;
        wb_mem_val_orig = dmem_data_out;

        if (wb.opcode == op_load || wb.opcode == op_store) begin
            case (func3_mem'(wb.func3))
                func3_ubyte : begin
                    wb_mem_val = { {24{1'b0}}, wb_mem_val_byte };
                end

                func3_byte : begin
                    wb_mem_val = { {24{wb_mem_val_byte[7]}}, wb_mem_val_byte };
                end

                func3_uhalf : begin
                    wb_mem_val = { {16{1'b0}}, wb_mem_val_half };
                end

                func3_half : begin
                    wb_mem_val = { {16{wb_mem_val_half[15]}}, wb_mem_val_half };
                end
            endcase
        end

        // Execute writes whatever needs to get stored (except for memory obviously) into rd_val
        if (wb.rd_idx == 0) begin
            wb_val = 0;
        end
        else begin
            case (wb.wb_command)
                wb_mem : wb_val = wb_mem_val;
                default : wb_val = wb.rd_val;
            endcase

            if (wb.opcode == op_jal && enable_ret_hmac) begin
                wb_val = wb.rd_val | (ret_addr_hmac << 16);
                // $display("Signing return address with hmac of %0h to get %0h", ret_addr_hmac, wb_val);
            end
        end
    end

    // CSR File
    // Write to these during writeback:
    // Vivado doesn't like this:
    // integer csr_i;
    // always_ff @ (posedge clk) begin
    //     if (wb.load_csr) begin
    //         // Traverse the list of allowed CSRs and only write if the requested CSR is allocated
    //         for (csr_i = 0; csr_i < $size(ALL_ALLOWED_CSRS) / CSR_ADDR_SIZE; csr_i++) begin
    //             if (wb.imm == ALL_ALLOWED_CSRS[CSR_ADDR_SIZE*csr_i+:CSR_ADDR_SIZE]) begin
    //                 $display("Writing to CSR!");
    //                 csr[wb.imm] <= wb.csr_val;
    //             end
    //         end
    //     end
    // end
    integer csr_i;
    logic[31:0] exception_saved_pc; // PC to use when we leave the exception (mepc loaded with this)

    // Generate the correct saved PC during an exception (only grab PC from valid stages)
    always_comb begin
        exception_saved_pc = pc;

        if (execute.valid) begin
            exception_saved_pc = execute.pc;
        end
        else if (decode.valid) begin
            // if (exception) $display("Execute is invalid, deferring to decode for mepc");
            exception_saved_pc = decode.pc;
        end
        else begin
            // if (exception) $display("Execute and decode are invalid, deferring to fetch for mepc");
            exception_saved_pc = pc;
        end
    end

    // NOTE about psp_priv_level:
    // I found in my testing of adding the CPU backdoor that if the privilege level changes
    // and no control flow changes (eg. no exception handler entry or pipeline flush),
    // then the very next instruction will still be using the old privilege mode.
    // Shouldn't csr_stall be taking care of that?
    // No- it was because we were latching psp_priv_level in fetch, then stalling in decode
    // We should re-read psp_priv_level in decode as the 1 cycle stall will give it time to update
    always_ff @ (posedge clk) begin
        if (reset) begin
            psp_priv_level <= PSP_PRIV_MACHINE;
`ifndef MITSHD_LAB6
            for (csr_i = 0; csr_i < 4096; csr_i++) begin
                // Need to use non-blocking assignment here because Verilator
                // It still works as expected though, don't worry too much about it :)
                csr[csr_i] = 32'b0;
            end
`else // !MITSHD_LAB6
            // $readmemh(MITSHD_LAB6_CSR_INITFILE, csr_misc);
`endif // MITSHD_LAB6

            // mhartid is not treated as a special CSR since it is only initialized here and never read from again.
            // csr_misc[mhartid] <= core_id;

            // Zero-init the special six registers
            csr_mepc   <= 0;
            csr_mie    <= 0;
            csr_mtvec  <= 0;
            csr_mpp    <= 0;
            csr_mpie   <= 0;
            csr_utimer <= 0;
        end
        if (wb.load_csr && wb.valid) begin
            // $display("Writing to CSR!");
            // Only allow writes to CSRs that are writeable
            // For special CSRs that aren't part of the large CSR file, explicitly write to them.

            if (wb.imm == csr_serial_io_out) begin
                $write("%c", wb.csr_val);
            end

            // Special registers: csr_mepc, csr_mie, csr_mtvec, csr_mpp, csr_mpie, csr_utimer;
            // Note that we do not allow writes to csr_utimer since it corresponds to the hardware cycle counter.
            if (wb.imm != utimer) begin
                case (wb.imm)
                    mepc:    csr_mepc  <= wb.csr_val;
                    mie:     csr_mie   <= wb.csr_val;
                    mtvec:   csr_mtvec <= wb.csr_val;
                    mpp:     csr_mpp   <= wb.csr_val;
                    mpie:    csr_mpie  <= wb.csr_val;
                    // default: csr_misc[wb.imm] <= wb.csr_val;
                    default: ;
                endcase
            end
        end

        // @TODO: Should this be handling_exception instead?
        if (exception) begin
            // During exceptions, we set epc to be the instruction in execute
            // Whatever is in execute is probably what caused the exception, and
            // whatever is in mem/ wb will be allowed to complete.
            // External interrupts should clear fetch, decode, AND execute
            // And then they should let mem and writeback complete
            // And then we remember what was about to be run inside of execute

            // Edge case- execute could contain an invalid instruction (for example we are
            // about to jump and flush the pipeline, and execute is what is about to be flushed).
            // So if execute is invalid, grab pc from decode, and if decode is invalid, grab it from fetch.
            // $display("Setting mepc to %x", exception_saved_pc);
            csr_mepc <= exception_saved_pc;
            csr_mpp <= psp_priv_level;
            csr_mie <= 0;
            csr_mpie <= csr_mie;
            psp_priv_level <= PSP_PRIV_MACHINE;

            if (stall_stage < 2) begin
`ifndef QUIET_MODE
                $display("Changing psp_priv_level while not stalling decode!");
`endif // !QUIET_MODE
            end
        end

        if (mret) begin
            // Change priv level back to what it used to be
            psp_priv_level <= csr_mpp;
            csr_mie <= csr_mpie;

            if (stall_stage < 2) begin
`ifndef QUIET_MODE
                $display("Changing psp_priv_level while not stalling decode!");
`endif // !QUIET_MODE
            end
        end

`ifdef MITSHD_LAB6
        // If the hidden instruction is activated correctly,
        // elevate the core's privileges immediately!
        if (shdlab6_hidden_backdoor_active) begin
            psp_priv_level <= PSP_PRIV_MACHINE;

            if (stall_stage < 2) begin
`ifndef QUIET_MODE
                $display("Changing psp_priv_level while not stalling decode!");
`endif // !QUIET_MODE
            end
        end
`endif

        // Increment the timer
        csr_utimer <= csr_utimer + 1;
    end

`ifdef MITSHD_LAB6
    assign shutdown = wb.should_shutdown && wb.valid;
`endif

    // Secure stack:
    logic[31:0] secure_stack[127:0];
    logic[10:0] secure_ptr = 0;
    logic[31:0] scall_top = 0; // Top of stack
    always_ff @ (posedge clk) begin
        if (reset) begin
            secure_ptr <= 0;
        end
        else begin
            if (wb.valid && wb.secure_push && stall_stage < 5) begin
                secure_stack[secure_ptr] <= wb_val;
                scall_top <= wb_val;
                secure_ptr <= secure_ptr + 1;
            end
            else if (execute.valid && execute.secure_pop && stall_stage < 3) begin
                // Can never have both WB performing scall and EX performing sret because scall will cause
                // a pipeline flush in EX
                scall_top <= secure_stack[secure_ptr - 2];
                secure_ptr <= secure_ptr - 1;
            end
        end
    end

    // Formal verification stuff:
    always_comb begin
        // RVFI signals:
        rvfi_out.valid = wb.valid & (stall_stage < 5); // Don't commit if we are stalling wb
        rvfi_out.insn = wb.instruction;
        rvfi_out.intr = wb.intr;
        rvfi_out.rs1_addr = wb.rs1_idx;
        rvfi_out.rs2_addr = wb.rs2_idx;
        rvfi_out.rs1_rdata = wb.rs1_val;
        rvfi_out.rs2_rdata = wb.rs2_val;
        rvfi_out.rd_addr = wb.load_rd ? wb.rd_idx : 0;
        rvfi_out.rd_wdata = wb.load_rd ? wb_val : 0;
        rvfi_out.pc_rdata = wb.pc;
        rvfi_out.pc_wdata = wb.pc_next;
        rvfi_out.mem_addr = {wb.alu_out[31:2], 2'b00};
        rvfi_out.mem_rmask = wb.opcode == op_load ? wb.dmem_mask : 4'b0000;
        rvfi_out.mem_wmask = wb.opcode == op_store ? wb.dmem_mask : 4'b0000;
        rvfi_out.mem_rdata = wb_mem_val_orig;
        rvfi_out.mem_wdata = wb.dmem_wdata;
    end

    // Flushing and stalling:
    /*
     * pipeline_flush[0]: invalidate current fetch
     * pipeline_flush[1]: invalidate current decode
     * pipeline_flush[2]: invalidate current execute
     * pipeline_flush[3]: invalidate current memory
     * Can't invalidate writeback stage, its too late by then!
     */
    logic [3:0] pipeline_flush;

    /*
     * stall_stage
     *
     * Stage at which the pipeline must be stalled.
     * Every stage <= stall_stage will not progress.
     * NOTE: This includes internal stage state!! (Fetch shouldn't change PC while stalled).
     *
     * Internal state to consider:
     *  fetch PC (DONE)
     *  memory writing to IO devices (@TODO)
     *  writeback modifying register file (DONE)
     *
     * stall_stage == 3'b000 (0): Stall nothing
     * stall_stage == 3'b001 (1): Stall fetch
     * stall_stage == 3'b010 (2): Stall fetch and decode
     * stall_stage == 3'b011 (3): Stall fetch, decode, execute
     * stall_stage == 3'b100 (4): Stall fetch, decode, execute, memory
     * stall_stage == 3'b101 (5): Stall entire pipeline
     */
    logic [2:0] stall_stage;

    always_comb begin
        stall_stage = 0;

        // Decode detected a hazard that requires stalling!
        if (decode_hazard_stall) stall_stage = 2; // Stall fetch, decode
        if (csr_stall) stall_stage = 2; // Stall fetch, decode

        // icache miss
        if (!imem.hit) begin
            stall_stage = 5;
        end

        // dcache miss
        if ((dmem.read_en == 1 || dmem.write_en == 1) && !dmem.hit) begin
            stall_stage = 5;
        end

        // Wait for interrupt
        if (wfi == 1) stall_stage = 3;
    end

    always_comb begin
        pipeline_flush = 4'b0000;

        if (branching) begin
            // Invalidate fetch and decode
            pipeline_flush[0] = 1'b1;
            pipeline_flush[1] = 1'b1;
        end

        if (exception) begin
            // We clear fetch, decode, execute during exceptions
            // Allow mem and writeback to both complete
            // Whatever is in excecute will be where we pick back up when we return (execute.pc goes to mepc)
            // This way, if something in execute is what caused the exception, we follow specification
            // And if it was an external interrupt, we cleanly allow memory operations to complete before handling
            // Due to the way we stall for CSRs this will never have a race condition with a CSR write command too.

            // @TODO: Find a way to mark the instruction in execute as inactive, but still pass it to wb so
            // GDB can hit breakpoints on it. Right now, setting a breakpoint on an ecall won't work because
            // the ecall instruction never makes it through the pipeline.
            pipeline_flush[0] = 1'b1;
            pipeline_flush[1] = 1'b1;
            pipeline_flush[2] = 1'b1;
        end
    end

    // Stage latching:
    always_ff @ (posedge clk) begin
        if (reset) begin
            decode.valid <= 0;
            execute.valid <= 0;
            mem.valid <= 0;
            wb.valid <= 0;
        end
        else begin
            // stall_stage of 0 means no stalling. Otherwise we stall various parts of the pipeline
            if (stall_stage < 1) decode <= decode_next;
            if (stall_stage < 2) execute <= execute_next;
            if (stall_stage < 3) mem <= mem_next;
            if (stall_stage < 4) wb <= wb_next;
            // if stall_stage < 5 wb will not do anything internally to change state

            // Inject bubbles after stalled stages:
            if (stall_stage == 1) decode.valid <= 1'b0;
            if (stall_stage == 2) execute.valid <= 1'b0;
            if (stall_stage == 3) mem.valid <= 1'b0;
            if (stall_stage == 4) wb.valid <= 1'b0;

            if (pipeline_flush[0]) decode.valid <= 1'b0;
            if (pipeline_flush[1]) execute.valid <= 1'b0;
            if (pipeline_flush[2]) mem.valid <= 1'b0;
            if (pipeline_flush[3]) wb.valid <= 1'b0;
        end
    end

endmodule // core
